*  Generated for: PrimeSim
*  Design library name: braun_mult
*  Design cell name: ks_adder_tb
*  Design view name: schematic
.lib 'saed32nm.lib' TT

*Custom Compiler Version S-2021.09
*Fri Feb 25 18:02:59 2022

.global gnd!
********************************************************************************
* Library          : braun_mult
* Cell             : cmosXOR
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosxor a_in b_in y_out
xm15 y_out net69 net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm7 net29 a_in net69 net29 p105 w=0.1u l=0.03u nf=1 m=1
xm6 net69 net13 net29 net29 p105 w=0.1u l=0.03u nf=1 m=1
xm5 net63 net50 net29 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm4 net29 b_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm2 net13 b_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm0 net50 a_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm16 y_out net69 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm11 gnd! a_in net44 gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm10 net47 net50 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm9 net44 net13 net69 net44 n105 w=0.1u l=0.03u nf=1 m=1
xm8 net69 b_in net47 net47 n105 w=0.1u l=0.03u nf=1 m=1
xm3 net13 b_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm1 net50 a_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
v17 net63 gnd! dc=1.8
.ends cmosxor

********************************************************************************
* Library          : braun_mult
* Cell             : cmosAND
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosand a_in b_in y_out
xm2 y_out net22 vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm1 net22 b_in vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm0 net22 a_in vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm5 net23 b_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm4 y_out net22 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm3 net22 a_in net23 net23 n105 w=0.1u l=0.03u nf=1 m=1
v9 vdd gnd! dc=1.8
.ends cmosand

********************************************************************************
* Library          : braun_mult
* Cell             : cmosOR
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosor a_in b_in out
xm4 out net25 net17 net17 p105 w=0.1u l=0.03u nf=1 m=1
xm2 net10 b_in net25 net10 p105 w=0.1u l=0.03u nf=1 m=1
xm1 net10 a_in net17 net17 p105 w=0.1u l=0.03u nf=1 m=1
xm6 net25 a_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm5 out net25 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm7 gnd! b_in net25 gnd! n105 w=0.1u l=0.03u nf=1 m=1
v8 net17 gnd! dc=1.8
.ends cmosor

********************************************************************************
* Library          : braun_mult
* Cell             : ks_adder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt ks_adder a0 a1 a2 b0 b1 b2 cin cout s0 s1 s2
xi21 net129 net116 s2 cmosxor
xi20 net130 net115 s1 cmosxor
xi19 cin net128 s0 cmosxor
xi12 a2 b2 net116 cmosxor
xi5 a1 b1 net115 cmosxor
xi0 a0 b0 net128 cmosxor
xi17 net121 net130 net76 cmosand
xi15 net115 net116 net121 cmosand
xi14 net116 net123 net125 cmosand
xi13 a2 b2 net127 cmosand
xi10 net120 cin net117 cmosand
xi8 net128 net115 net120 cmosand
xi7 net115 net122 net126 cmosand
xi6 a1 b1 net123 cmosand
xi2 cin net128 net124 cmosand
xi1 a0 b0 net122 cmosand
xi18 net76 net119 cout cmosor
xi16 net125 net127 net119 cmosor
xi11 net117 net118 net129 cmosor
xi9 net126 net123 net118 cmosor
xi3 net124 net122 net130 cmosor
.ends ks_adder

********************************************************************************
* Library          : braun_mult
* Cell             : ks_adder_tb
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
xi0 a0 a1 a2 b0 b1 b2 cin cout s0 s1 s2 ks_adder
v7 a0 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 5u 10u )
v6 a1 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 10u 20u )
v5 a2 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 15u 30u )
v4 b0 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 20u 40u )
v3 b1 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 25u 50u )
v2 b2 gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 30u 60u )
v1 cin gnd! dc=0 pulse ( 1.8 0 0 0.1n 0.1n 35u 70u )








.tran '0.1u' '140u' name=tran

.option primesim_remove_probe_prefix = 0
.probe v(*) i(*) level=1
.probe tran v(a0) v(a1) v(a2) v(b0) v(b1) v(b2) v(cin) v(cout) v(s0) v(s1) v(s2)

.temp 25



.option primesim_output=wdf


.option parhier = LOCAL






.end
