*  Generated for: PrimeSim
*  Design library name: braun_mult
*  Design cell name: braun_multiplier_tb
*  Design view name: schematic
.lib 'saed32nm.lib' TT

*Custom Compiler Version S-2021.09
*Fri Feb 25 18:33:07 2022

.global gnd!
********************************************************************************
* Library          : braun_mult
* Cell             : cmosAND
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosand a_in b_in y_out
xm2 y_out net22 vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm1 net22 b_in vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm0 net22 a_in vdd vdd p105 w=0.1u l=0.03u nf=1 m=1
xm5 net23 b_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm4 y_out net22 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm3 net22 a_in net23 net23 n105 w=0.1u l=0.03u nf=1 m=1
v9 vdd gnd! dc=1.8
.ends cmosand

********************************************************************************
* Library          : braun_mult
* Cell             : cmosXOR
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosxor a_in b_in y_out
xm15 y_out net69 net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm7 net29 a_in net69 net29 p105 w=0.1u l=0.03u nf=1 m=1
xm6 net69 net13 net29 net29 p105 w=0.1u l=0.03u nf=1 m=1
xm5 net63 net50 net29 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm4 net29 b_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm2 net13 b_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm0 net50 a_in net63 net63 p105 w=0.1u l=0.03u nf=1 m=1
xm16 y_out net69 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm11 gnd! a_in net44 gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm10 net47 net50 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm9 net44 net13 net69 net44 n105 w=0.1u l=0.03u nf=1 m=1
xm8 net69 b_in net47 net47 n105 w=0.1u l=0.03u nf=1 m=1
xm3 net13 b_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm1 net50 a_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
v17 net63 gnd! dc=1.8
.ends cmosxor

********************************************************************************
* Library          : braun_mult
* Cell             : half_adder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt half_adder carry sum x y
xi0 x y sum cmosxor
xi1 x y carry cmosand
.ends half_adder

********************************************************************************
* Library          : braun_mult
* Cell             : full_adder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt full_adder c_in carry sum x_in y_in
xi1 net20 sum net22 c_in half_adder
xi0 net21 net22 x_in y_in half_adder
xi2 net21 net20 carry cmosxor
.ends full_adder

********************************************************************************
* Library          : braun_mult
* Cell             : cmosOR
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt cmosor a_in b_in out
xm4 out net25 net17 net17 p105 w=0.1u l=0.03u nf=1 m=1
xm2 net10 b_in net25 net10 p105 w=0.1u l=0.03u nf=1 m=1
xm1 net10 a_in net17 net17 p105 w=0.1u l=0.03u nf=1 m=1
xm6 net25 a_in gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm5 out net25 gnd! gnd! n105 w=0.1u l=0.03u nf=1 m=1
xm7 gnd! b_in net25 gnd! n105 w=0.1u l=0.03u nf=1 m=1
v8 net17 gnd! dc=1.8
.ends cmosor

********************************************************************************
* Library          : braun_mult
* Cell             : ks_adder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt ks_adder a0 a1 a2 b0 b1 b2 cin cout s0 s1 s2
xi21 net129 net116 s2 cmosxor
xi20 net130 net115 s1 cmosxor
xi19 cin net128 s0 cmosxor
xi12 a2 b2 net116 cmosxor
xi5 a1 b1 net115 cmosxor
xi0 a0 b0 net128 cmosxor
xi17 net121 net130 net76 cmosand
xi15 net115 net116 net121 cmosand
xi14 net116 net123 net125 cmosand
xi13 a2 b2 net127 cmosand
xi10 net120 cin net117 cmosand
xi8 net128 net115 net120 cmosand
xi7 net115 net122 net126 cmosand
xi6 a1 b1 net123 cmosand
xi2 cin net128 net124 cmosand
xi1 a0 b0 net122 cmosand
xi18 net76 net119 cout cmosor
xi16 net125 net127 net119 cmosor
xi11 net117 net118 net129 cmosor
xi9 net126 net123 net118 cmosor
xi3 net124 net122 net130 cmosor
.ends ks_adder

********************************************************************************
* Library          : braun_mult
* Cell             : braun_multiplier
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt braun_multiplier p0 p1 p2 p3 p4 p5 p6 p7 x0 x1 x2 x3 y0 y1 y2 y3
xi32 x0 y3 net174 cmosand
xi31 x1 y3 net170 cmosand
xi30 x2 y3 net81 cmosand
xi5 x2 y1 net156 cmosand
xi18 x3 y3 net105 cmosand
xi14 x0 y2 net166 cmosand
xi13 x1 y2 net164 cmosand
xi12 x2 y2 net162 cmosand
xi11 x3 y2 net83 cmosand
xi7 x0 y1 net160 cmosand
xi6 x1 y1 net158 cmosand
xi4 x3 y1 net56 cmosand
xi3 x0 y0 p0 cmosand
xi2 x1 y0 net39 cmosand
xi1 x2 y0 net34 cmosand
xi0 x3 y0 net29 cmosand
xi24 net89 net96 p3 net174 net93 full_adder
xi23 net84 net97 net101 net170 net88 full_adder
xi22 net79 net99 net103 net81 net83 full_adder
xi17 net62 net89 p2 net166 net94 full_adder
xi16 net57 net84 net93 net164 net61 full_adder
xi15 net52 net79 net88 net162 net56 full_adder
xi10 gnd! net62 p1 net160 net39 full_adder
xi9 gnd! net57 net94 net158 net34 full_adder
xi8 gnd! net52 net61 net156 net29 full_adder
xi25 net96 net97 net99 net101 net103 net105 gnd! p7 p4 p5 p6 ks_adder
.ends braun_multiplier

********************************************************************************
* Library          : braun_mult
* Cell             : braun_multiplier_tb
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
xi0 p0 p1 p2 p3 p4 p5 p6 p7 x0 x1 x2 x3 y0 y1 y2 y3 braun_multiplier
v8 y3 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 5u 10u )
v7 y2 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 40u 80u )
v6 y1 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 20u 40u )
v5 y0 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 10u 20u )
v4 x3 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 5u 10u )
v3 x2 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 10u 20u )
v2 x1 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 20u 40u )
v1 x0 gnd! dc=0 pulse ( 0 1.8 0 0.1n 0.1n 40u 80u )








.tran '0.1u' '100u' name=tran

.option primesim_remove_probe_prefix = 0
.probe v(*) i(*) level=1
.probe tran v(x0) v(x1) v(x2) v(x3) v(y0) v(y1) v(y2) v(y3) v(p0) v(p1) v(p2) v(p3) v(p4) v(p5) v(p6) v(p7)

.temp 25



.option primesim_output=wdf


.option parhier = LOCAL






.end
